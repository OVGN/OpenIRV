/* 
 * ----------------------------------------------------------------------------
 *  Project:  OpenIRV
 *  Filename: i2c_eeprom_emulator.v
 *  Purpose:  Current module allows to emulate I2C EEPROM. 
 * ----------------------------------------------------------------------------
 *  Copyright © 2020-2021, Vaagn Oganesyan <ovgn@protonmail.com>
 *  
 *  Licensed under the Apache License, Version 2.0 (the "License");
 *  you may not use this file except in compliance with the License.
 *  You may obtain a copy of the License at
 *  
 *      http://www.apache.org/licenses/LICENSE-2.0
 *  
 *  Unless required by applicable law or agreed to in writing, software
 *  distributed under the License is distributed on an "AS IS" BASIS,
 *  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *  See the License for the specific language governing permissions and
 * ----------------------------------------------------------------------------
 */


`default_nettype none
`timescale 1ps / 1ps


module i2c_eeprom_emulator #
(
    parameter   [6:0]   EEPROM_I2C_ADDRESS = 7'b1010001,
    parameter           WR_ENA = 1'b1
)
(
    input   wire    clk,
    input   wire    rstn,

    (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME LUT_RAM, MEM_SIZE 4096, MASTER_TYPE BRAM_CTRL, MEM_WIDTH 32, MEM_ECC NONE, READ_LATENCY 1, READ_WRITE_MODE READ_WRITE" *)
    (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 EMU_RAM CLK"   *)  input   wire            bram_clk,
    (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 EMU_RAM EN "   *)  input   wire            bram_ena,
    (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 EMU_RAM RST"   *)  input   wire            bram_rst,
    (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 EMU_RAM WE"    *)  input   wire    [3:0]   bram_we,
    (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 EMU_RAM ADDR"  *)  input   wire    [31:0]  bram_addr,
    (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 EMU_RAM DIN"   *)  input   wire    [31:0]  bram_wdata,
    (* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 EMU_RAM DOUT"  *)  output  wire    [31:0]  bram_rdata,

    (* X_INTERFACE_INFO = "xilinx.com:interface:iic:1.0 IIC SCL_I" *)       input   wire    scl_i,
    (* X_INTERFACE_INFO = "xilinx.com:interface:iic:1.0 IIC SCL_O" *)       output  wire    scl_o,
    (* X_INTERFACE_INFO = "xilinx.com:interface:iic:1.0 IIC SCL_T" *)       output  wire    scl_t,
    (* X_INTERFACE_INFO = "xilinx.com:interface:iic:1.0 IIC SDA_I" *)       input   wire    sda_i,
    (* X_INTERFACE_INFO = "xilinx.com:interface:iic:1.0 IIC SDA_O" *)       output  wire    sda_o,
    (* X_INTERFACE_INFO = "xilinx.com:interface:iic:1.0 IIC SDA_T" *)       output  reg     sda_t = 1'b1
);

/*-------------------------------------------------------------------------------------------------------------------------------------*/
    
    wire scl;
    wire sda;
    
    sync_cdc_bit #
    (
        .C_SYNC_STAGES (3)
    )
    sync_cdc_bit_scl
    (
        .clk ( clk   ),
        .d   ( scl_i ),
        .q   ( scl   )
    );
    
    
    sync_cdc_bit #
    (
        .C_SYNC_STAGES (3)
    )
    sync_cdc_bit_sda
    (
        .clk ( clk   ),
        .d   ( sda_i ),
        .q   ( sda   )
    );

/*-------------------------------------------------------------------------------------------------------------------------------------*/
    
    reg     scl_1 = 1'b1;
    reg     sda_1 = 1'b1;
    
    reg     scl_fe = 1'b0;
    reg     sda_fe = 1'b0;
    
    reg     scl_re = 1'b0;
    reg     sda_re = 1'b0;
    
    reg     i2c_start = 1'b0;
    reg     i2c_stop  = 1'b0;
    
    
    always @(posedge clk) begin
        if (~rstn) begin
            scl_1     <= 1'b1;
            sda_1     <= 1'b1;
            scl_fe    <= 1'b0;
            sda_fe    <= 1'b0;
            scl_re    <= 1'b0;
            sda_re    <= 1'b0;
            i2c_start <= 1'b0;
            i2c_stop  <= 1'b0;
        end else begin
            scl_1 <= scl;
            sda_1 <= sda;
            
            scl_fe <=  scl_1 & ~scl;
            scl_re <= ~scl_1 &  scl;
            
            sda_fe <=  sda_1 & ~sda;
            sda_re <= ~sda_1 &  sda;
            
            i2c_start <= sda_fe & scl;
            i2c_stop  <= sda_re & scl;
        end
    end

/*-------------------------------------------------------------------------------------------------------------------------------------*/
    
    wire    scl_fe_delayed;
    
    /* Current delay after SCL falling edge
     * allows to prevent false START bus 
     * condition generated by slave device */
    pipeline #
    (
        .PIPE_WIDTH ( 1  ),
        .PIPE_STAGES( 10 )      // TODO: this value depends on the system to I2C clock speed ratio
    )
    pipeline_inst
    (
        .clk        ( clk            ), 
        .cen        ( 1'b1           ), 
        .srst       ( ~rstn          ), 
        .pipe_in    ( scl_fe         ), 
        .pipe_out   ( scl_fe_delayed )
    );

/*-------------------------------------------------------------------------------------------------------------------------------------*/
    
    reg     [7:0]   cnt  = 8'h00;
    reg     [7:0]   din  = 8'h00;
    reg     [7:0]   dout = 8'h00;
    reg     [7:0]   mem_addr_high = 8'h00;
    reg     [7:0]   mem_addr_low  = 8'h00;
    
    reg             ram_we   = 1'b0;
    reg     [15:0]  ram_addr = 16'h0000;
    reg     [7:0]   ram_din  = 8'h00;
    wire    [7:0]   ram_dout;
    
    
    localparam  [2:0]   ST_STOP             = 3'd0,
                        ST_START            = 3'd1,
                        ST_CHECK_SLAVE_ADDR = 3'd2,
                        ST_SEND_ACK         = 3'd3,
                        ST_MEM_ADDR_HIGH    = 3'd4,
                        ST_MEM_ADDR_LOW     = 3'd5,
                        ST_MEM_READ         = 3'd6,
                        ST_MEM_WRITE        = 3'd7;
    
    reg     [2:0]   state      = ST_STOP;
    reg     [2:0]   next_state = ST_STOP;
    
    
    always @(posedge clk) begin
        if (~rstn) begin
            ram_we <= 1'b0;
            sda_t  <= 1'b1;
            state  <= ST_STOP;
        end else begin
            
            /* Start and stop bus conditions have higher
             * priority over all other states and events */
            if (i2c_start) begin
                state <= ST_START;
            end else begin
                if (i2c_stop) begin
                    state <= ST_STOP;
                end else begin
                    case (state)
                        
                        ST_STOP: begin
                            sda_t <= 1'b1;
                            state <= state;
                        end
                        
                        ST_START: begin
                            sda_t <= 1'b1;
                            cnt   <= 8'd0;
                            state <= ST_CHECK_SLAVE_ADDR;
                        end
                        
                        ST_CHECK_SLAVE_ADDR: begin
                            if (cnt < 8'd8) begin
                                if (scl_re) begin
                                    cnt <= cnt + 1'b1;
                                    din <= {din[6:0], sda};
                                end
                            end else begin
                                if (din[7:1] == EEPROM_I2C_ADDRESS) begin
                                    if (scl_fe_delayed) begin
                                        sda_t <= ram_dout[7];
                                        dout  <= {ram_dout[6:0], ram_dout[7]};
                                        state <= ST_SEND_ACK;
                                        next_state <= (din[0])? ST_MEM_READ : ST_MEM_ADDR_HIGH;
                                    end
                                end else begin
                                    state <= ST_STOP;
                                end
                            end
                        end
                        
                        ST_SEND_ACK: begin
                            cnt <= 8'd0;
                            if (scl_fe_delayed) begin
                                state <= next_state;
                                sda_t <= 1'b1;
                            end else begin
                                sda_t <= 1'b0;
                            end
                        end
                        
                        ST_MEM_ADDR_HIGH: begin
                            if (cnt < 8'd8) begin
                                if (scl_re) begin
                                    cnt <= cnt + 1'b1;
                                    mem_addr_high <= {mem_addr_high[6:0], sda};
                                end
                            end else begin
                                if (scl_fe_delayed) begin
                                    state <= ST_SEND_ACK;
                                    next_state <= ST_MEM_ADDR_LOW;
                                end
                            end
                        end
                        
                        ST_MEM_ADDR_LOW: begin
                            if (cnt < 8'd8) begin
                                if (scl_re) begin
                                    cnt <= cnt + 1'b1;
                                    mem_addr_low <= {mem_addr_low[6:0], sda};
                                end
                            end else begin
                                if (scl_fe_delayed) begin
                                    ram_addr <= {mem_addr_high, mem_addr_low};
                                    state <= ST_SEND_ACK;
                                    next_state <= ST_MEM_WRITE;
                                end
                            end
                        end
                        
                        ST_MEM_READ: begin
                            if (cnt < 8'd8) begin
                                if (cnt < 8'd7) begin
                                    if (scl_fe_delayed) begin
                                        sda_t <= dout[7];
                                        cnt <= cnt + 1'b1;
                                        dout <= {dout[6:0], dout[7]};
                                    end
                                end else begin
                                    /* Stop driving SDA line, to get ACK from master */
                                    if (scl_fe_delayed) begin
                                        cnt <= cnt + 1'b1;
                                        sda_t <= 1'b1;
                                    end
                                end
                            end else begin
                                /* Check ACK from master to continue or stop reading */
                                if (scl_re) begin
                                    ram_addr <= ram_addr + 1'b1;
                                    next_state <= (sda)? ST_STOP : ST_MEM_READ;
                                end
                                
                                if (scl_fe_delayed) begin
                                    cnt <= 8'd0;
                                    sda_t <= ram_dout[7];
                                    dout  <= {ram_dout[6:0], ram_dout[7]};
                                    state <= next_state;
                                end
                            end
                        end
                        
                        ST_MEM_WRITE: begin
                            if (cnt < 8'd8) begin
                                if (scl_re) begin
                                    cnt <= cnt + 1'b1;
                                    ram_din <= {ram_din[6:0], sda};
                                end
                            end else begin
                                if (scl_fe_delayed) begin
                                    ram_we <= 1'b1;
                                end
                                
                                if (ram_we) begin
                                    ram_we <= 1'b0;
                                    ram_addr <= ram_addr + 1'b1;
                                    state <= ST_SEND_ACK;
                                    next_state <= ST_MEM_WRITE;
                                end
                            end
                        end
                        
                        default: begin
                            state <= ST_STOP;
                        end
                        
                    endcase
                end
            end
        end
    end
    
/*-------------------------------------------------------------------------------------------------------------------------------------*/
    
    I2C_EEPROM_EMU_RAM I2C_EEPROM_EMU_RAM_inst
    (
        .clka   ( bram_clk        ),    // input wire clka
        .rsta   ( bram_rst        ),    // input wire rsta
        .ena    ( bram_ena        ),    // input wire ena
        .wea    ( bram_we         ),    // input wire [3 : 0] wea
        .addra  ( bram_addr[11:2] ),    // input wire [9 : 0] addra
        .dina   ( bram_wdata      ),    // input wire [31 : 0] dina
        .douta  ( bram_rdata      ),    // output wire [31 : 0] douta
        
        .clkb   ( clk             ),    // input wire clkb
        .rstb   ( 1'b0            ),    // input wire rstb
        .enb    ( 1'b1            ),    // input wire enb
        .web    ( ram_we & WR_ENA ),    // input wire [0 : 0] web
        .addrb  ( ram_addr[11:0]  ),    // input wire [11 : 0] addrb
        .dinb   ( ram_din         ),    // input wire [7 : 0] dinb
        .doutb  ( ram_dout        )     // output wire [7 : 0] doutb
    );
    
/*-------------------------------------------------------------------------------------------------------------------------------------*/
    
    assign scl_o = 1'b0;
    assign scl_t = 1'b1;
    assign sda_o = 1'b0;
    
endmodule

/*-------------------------------------------------------------------------------------------------------------------------------------*/

`default_nettype wire
